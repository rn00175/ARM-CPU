module prog_counter ()